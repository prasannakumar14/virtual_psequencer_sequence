package pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;
 
  `include "xtn.sv"
  `include "agent_config.sv"
  `include "sequencer.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "agent.sv"
  `include "seqs.sv"
  `include "virtual_sequencer.sv"
  `include "virtual_sequence.sv"

  `include "env.sv"
  `include "test.sv"
endpackage

